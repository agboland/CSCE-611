/* Control Unit implementation */
module ControlUnit (
    input wire 
    input wire [11:0] address,
    output wire [31:0] instruction
);